// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		inout  wire        av_config_SDAT,                          //                        av_config.SDAT
		output wire        av_config_SCLK,                          //                                 .SCLK
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,         //                           hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,           //                                 .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,           //                                 .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,           //                                 .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,           //                                 .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,           //                                 .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,           //                                 .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,            //                                 .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,         //                                 .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,         //                                 .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,         //                                 .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,           //                                 .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,           //                                 .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,           //                                 .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,             //                                 .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,             //                                 .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,             //                                 .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,             //                                 .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,             //                                 .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,             //                                 .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,             //                                 .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,              //                                 .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,              //                                 .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,             //                                 .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,              //                                 .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,              //                                 .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,              //                                 .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,              //                                 .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,              //                                 .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,              //                                 .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,              //                                 .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,              //                                 .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,              //                                 .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,              //                                 .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,             //                                 .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,             //                                 .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,             //                                 .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,             //                                 .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,            //                                 .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,           //                                 .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,           //                                 .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,            //                                 .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,             //                                 .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,             //                                 .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,             //                                 .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,             //                                 .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,             //                                 .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,             //                                 .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,          //                                 .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,          //                                 .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,          //                                 .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,          //                                 .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,          //                                 .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,          //                                 .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,          //                                 .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,          //                                 .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                            //                           memory.mem_a
		output wire [2:0]  memory_mem_ba,                           //                                 .mem_ba
		output wire        memory_mem_ck,                           //                                 .mem_ck
		output wire        memory_mem_ck_n,                         //                                 .mem_ck_n
		output wire        memory_mem_cke,                          //                                 .mem_cke
		output wire        memory_mem_cs_n,                         //                                 .mem_cs_n
		output wire        memory_mem_ras_n,                        //                                 .mem_ras_n
		output wire        memory_mem_cas_n,                        //                                 .mem_cas_n
		output wire        memory_mem_we_n,                         //                                 .mem_we_n
		output wire        memory_mem_reset_n,                      //                                 .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                           //                                 .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                          //                                 .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                        //                                 .mem_dqs_n
		output wire        memory_mem_odt,                          //                                 .mem_odt
		output wire [3:0]  memory_mem_dm,                           //                                 .mem_dm
		input  wire        memory_oct_rzqin,                        //                                 .oct_rzqin
		output wire [12:0] sdram_addr,                              //                            sdram.addr
		output wire [1:0]  sdram_ba,                                //                                 .ba
		output wire        sdram_cas_n,                             //                                 .cas_n
		output wire        sdram_cke,                               //                                 .cke
		output wire        sdram_cs_n,                              //                                 .cs_n
		inout  wire [15:0] sdram_dq,                                //                                 .dq
		output wire [1:0]  sdram_dqm,                               //                                 .dqm
		output wire        sdram_ras_n,                             //                                 .ras_n
		output wire        sdram_we_n,                              //                                 .we_n
		output wire        sdram_clk_clk,                           //                        sdram_clk.clk
		input  wire        system_pll_ref_clk_clk,                  //               system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,              //             system_pll_ref_reset.reset
		output wire        vga_CLK,                                 //                              vga.CLK
		output wire        vga_HS,                                  //                                 .HS
		output wire        vga_VS,                                  //                                 .VS
		output wire        vga_BLANK,                               //                                 .BLANK
		output wire        vga_SYNC,                                //                                 .SYNC
		output wire [7:0]  vga_R,                                   //                                 .R
		output wire [7:0]  vga_G,                                   //                                 .G
		output wire [7:0]  vga_B,                                   //                                 .B
		input  wire        vga_pll_ref_clk_clk,                     //                  vga_pll_ref_clk.clk
		input  wire        vga_pll_ref_reset_reset,                 //                vga_pll_ref_reset.reset
		output wire [31:0] x_coordinate_external_connection_export, // x_coordinate_external_connection.export
		output wire [31:0] y_coordinate_external_connection_export  // y_coordinate_external_connection.export
	);

	wire          system_pll_sys_clk_clk;                                               // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, AV_Config:clk, Onchip_SRAM:clk, Pixel_DMA_Addr_Translation:clk, SDRAM:clk, VGA_Subsystem:sys_clk_clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, mm_interconnect_2:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_002:clk, x_coordinate:clk, y_coordinate:clk]
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;                                    // ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;                                      // ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;                                      // ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_wready;                                     // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;                                        // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_rready;                                     // ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;                                      // ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;                                        // ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;                                    // ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	wire          arm_a9_hps_h2f_axi_master_wvalid;                                     // ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;                                     // ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;                                     // ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;                                     // ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;                                      // ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_arvalid;                                    // ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;                                    // ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;                                       // ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;                                     // ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;                                     // ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;                                     // ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	wire          arm_a9_hps_h2f_axi_master_arready;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	wire          arm_a9_hps_h2f_axi_master_awready;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;                                    // ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;                                     // ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	wire          arm_a9_hps_h2f_axi_master_bready;                                     // ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	wire          arm_a9_hps_h2f_axi_master_rlast;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	wire          arm_a9_hps_h2f_axi_master_wlast;                                      // ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;                                       // ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;                                        // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	wire          arm_a9_hps_h2f_axi_master_bvalid;                                     // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;                                     // ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	wire          arm_a9_hps_h2f_axi_master_awvalid;                                    // ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	wire          arm_a9_hps_h2f_axi_master_rvalid;                                     // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	wire          vga_subsystem_pixel_dma_master_waitrequest;                           // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	wire   [15:0] vga_subsystem_pixel_dma_master_readdata;                              // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	wire   [31:0] vga_subsystem_pixel_dma_master_address;                               // VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_address
	wire          vga_subsystem_pixel_dma_master_read;                                  // VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_read
	wire          vga_subsystem_pixel_dma_master_readdatavalid;                         // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	wire          vga_subsystem_pixel_dma_master_lock;                                  // VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_lock
	wire          mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect;         // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_chipselect -> VGA_Subsystem:char_buffer_slave_chipselect
	wire    [7:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata;           // VGA_Subsystem:char_buffer_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_slave_readdata
	wire          mm_interconnect_0_vga_subsystem_char_buffer_slave_waitrequest;        // VGA_Subsystem:char_buffer_slave_waitrequest -> mm_interconnect_0:VGA_Subsystem_char_buffer_slave_waitrequest
	wire   [12:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_address;            // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_address -> VGA_Subsystem:char_buffer_slave_address
	wire          mm_interconnect_0_vga_subsystem_char_buffer_slave_read;               // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_read -> VGA_Subsystem:char_buffer_slave_read
	wire    [0:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable;         // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_byteenable -> VGA_Subsystem:char_buffer_slave_byteenable
	wire          mm_interconnect_0_vga_subsystem_char_buffer_slave_write;              // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_write -> VGA_Subsystem:char_buffer_slave_write
	wire    [7:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata;          // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_writedata -> VGA_Subsystem:char_buffer_slave_writedata
	wire          mm_interconnect_0_sdram_s1_chipselect;                                // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire   [15:0] mm_interconnect_0_sdram_s1_readdata;                                  // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire          mm_interconnect_0_sdram_s1_waitrequest;                               // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire   [24:0] mm_interconnect_0_sdram_s1_address;                                   // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire          mm_interconnect_0_sdram_s1_read;                                      // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire    [1:0] mm_interconnect_0_sdram_s1_byteenable;                                // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire          mm_interconnect_0_sdram_s1_readdatavalid;                             // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire          mm_interconnect_0_sdram_s1_write;                                     // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire   [15:0] mm_interconnect_0_sdram_s1_writedata;                                 // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire          mm_interconnect_0_onchip_sram_s2_chipselect;                          // mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	wire    [7:0] mm_interconnect_0_onchip_sram_s2_readdata;                            // Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	wire   [16:0] mm_interconnect_0_onchip_sram_s2_address;                             // mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	wire          mm_interconnect_0_onchip_sram_s2_write;                               // mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	wire    [7:0] mm_interconnect_0_onchip_sram_s2_writedata;                           // mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	wire          mm_interconnect_0_onchip_sram_s2_clken;                               // mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                                 // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                   // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                   // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire          arm_a9_hps_h2f_lw_axi_master_wready;                                  // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                     // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire          arm_a9_hps_h2f_lw_axi_master_rready;                                  // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                   // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                     // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                                 // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire          arm_a9_hps_h2f_lw_axi_master_wvalid;                                  // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                  // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                  // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                  // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                   // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire          arm_a9_hps_h2f_lw_axi_master_arvalid;                                 // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                                 // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                    // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                  // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                  // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                  // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                   // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire          arm_a9_hps_h2f_lw_axi_master_arready;                                 // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                   // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire          arm_a9_hps_h2f_lw_axi_master_awready;                                 // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                                 // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                  // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire          arm_a9_hps_h2f_lw_axi_master_bready;                                  // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire          arm_a9_hps_h2f_lw_axi_master_rlast;                                   // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire          arm_a9_hps_h2f_lw_axi_master_wlast;                                   // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                   // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                    // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                     // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire          arm_a9_hps_h2f_lw_axi_master_bvalid;                                  // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                  // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire          arm_a9_hps_h2f_lw_axi_master_awvalid;                                 // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire          arm_a9_hps_h2f_lw_axi_master_rvalid;                                  // mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_av_config_avalon_av_config_slave_readdata;          // AV_Config:readdata -> mm_interconnect_1:AV_Config_avalon_av_config_slave_readdata
	wire          mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest;       // AV_Config:waitrequest -> mm_interconnect_1:AV_Config_avalon_av_config_slave_waitrequest
	wire    [1:0] mm_interconnect_1_av_config_avalon_av_config_slave_address;           // mm_interconnect_1:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire          mm_interconnect_1_av_config_avalon_av_config_slave_read;              // mm_interconnect_1:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire    [3:0] mm_interconnect_1_av_config_avalon_av_config_slave_byteenable;        // mm_interconnect_1:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire          mm_interconnect_1_av_config_avalon_av_config_slave_write;             // mm_interconnect_1:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire   [31:0] mm_interconnect_1_av_config_avalon_av_config_slave_writedata;         // mm_interconnect_1:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire          mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect; // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_chipselect -> VGA_Subsystem:char_buffer_control_slave_chipselect
	wire   [31:0] mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata;   // VGA_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_readdata
	wire    [0:0] mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address;    // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_address -> VGA_Subsystem:char_buffer_control_slave_address
	wire          mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read;       // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_read -> VGA_Subsystem:char_buffer_control_slave_read
	wire    [3:0] mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable; // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_byteenable -> VGA_Subsystem:char_buffer_control_slave_byteenable
	wire          mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write;      // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_write -> VGA_Subsystem:char_buffer_control_slave_write
	wire   [31:0] mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata;  // mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_writedata -> VGA_Subsystem:char_buffer_control_slave_writedata
	wire          mm_interconnect_1_x_coordinate_s1_chipselect;                         // mm_interconnect_1:x_coordinate_s1_chipselect -> x_coordinate:chipselect
	wire   [31:0] mm_interconnect_1_x_coordinate_s1_readdata;                           // x_coordinate:readdata -> mm_interconnect_1:x_coordinate_s1_readdata
	wire    [1:0] mm_interconnect_1_x_coordinate_s1_address;                            // mm_interconnect_1:x_coordinate_s1_address -> x_coordinate:address
	wire          mm_interconnect_1_x_coordinate_s1_write;                              // mm_interconnect_1:x_coordinate_s1_write -> x_coordinate:write_n
	wire   [31:0] mm_interconnect_1_x_coordinate_s1_writedata;                          // mm_interconnect_1:x_coordinate_s1_writedata -> x_coordinate:writedata
	wire          mm_interconnect_1_y_coordinate_s1_chipselect;                         // mm_interconnect_1:y_coordinate_s1_chipselect -> y_coordinate:chipselect
	wire   [31:0] mm_interconnect_1_y_coordinate_s1_readdata;                           // y_coordinate:readdata -> mm_interconnect_1:y_coordinate_s1_readdata
	wire    [1:0] mm_interconnect_1_y_coordinate_s1_address;                            // mm_interconnect_1:y_coordinate_s1_address -> y_coordinate:address
	wire          mm_interconnect_1_y_coordinate_s1_write;                              // mm_interconnect_1:y_coordinate_s1_write -> y_coordinate:write_n
	wire   [31:0] mm_interconnect_1_y_coordinate_s1_writedata;                          // mm_interconnect_1:y_coordinate_s1_writedata -> y_coordinate:writedata
	wire   [31:0] mm_interconnect_1_pixel_dma_addr_translation_slave_readdata;          // Pixel_DMA_Addr_Translation:slave_readdata -> mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_readdata
	wire          mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest;       // Pixel_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_waitrequest
	wire    [1:0] mm_interconnect_1_pixel_dma_addr_translation_slave_address;           // mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_address -> Pixel_DMA_Addr_Translation:slave_address
	wire          mm_interconnect_1_pixel_dma_addr_translation_slave_read;              // mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_read -> Pixel_DMA_Addr_Translation:slave_read
	wire    [3:0] mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable;        // mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_byteenable -> Pixel_DMA_Addr_Translation:slave_byteenable
	wire          mm_interconnect_1_pixel_dma_addr_translation_slave_write;             // mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_write -> Pixel_DMA_Addr_Translation:slave_write
	wire   [31:0] mm_interconnect_1_pixel_dma_addr_translation_slave_writedata;         // mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_writedata -> Pixel_DMA_Addr_Translation:slave_writedata
	wire   [31:0] pixel_dma_addr_translation_master_readdata;                           // mm_interconnect_2:Pixel_DMA_Addr_Translation_master_readdata -> Pixel_DMA_Addr_Translation:master_readdata
	wire          pixel_dma_addr_translation_master_waitrequest;                        // mm_interconnect_2:Pixel_DMA_Addr_Translation_master_waitrequest -> Pixel_DMA_Addr_Translation:master_waitrequest
	wire    [1:0] pixel_dma_addr_translation_master_address;                            // Pixel_DMA_Addr_Translation:master_address -> mm_interconnect_2:Pixel_DMA_Addr_Translation_master_address
	wire    [3:0] pixel_dma_addr_translation_master_byteenable;                         // Pixel_DMA_Addr_Translation:master_byteenable -> mm_interconnect_2:Pixel_DMA_Addr_Translation_master_byteenable
	wire          pixel_dma_addr_translation_master_read;                               // Pixel_DMA_Addr_Translation:master_read -> mm_interconnect_2:Pixel_DMA_Addr_Translation_master_read
	wire          pixel_dma_addr_translation_master_write;                              // Pixel_DMA_Addr_Translation:master_write -> mm_interconnect_2:Pixel_DMA_Addr_Translation_master_write
	wire   [31:0] pixel_dma_addr_translation_master_writedata;                          // Pixel_DMA_Addr_Translation:master_writedata -> mm_interconnect_2:Pixel_DMA_Addr_Translation_master_writedata
	wire   [31:0] mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_readdata;     // VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_address;      // mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	wire          mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_read;         // mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	wire    [3:0] mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_byteenable;   // mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	wire          mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_write;        // mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	wire   [31:0] mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_writedata;    // mm_interconnect_2:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                                              // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                                              // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [AV_Config:reset, Onchip_SRAM:reset, Pixel_DMA_Addr_Translation:reset, SDRAM:reset_n, mm_interconnect_0:SDRAM_reset_reset_bridge_in_reset_reset, mm_interconnect_0:VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:AV_Config_reset_reset_bridge_in_reset_reset, mm_interconnect_1:VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_2:Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset, mm_interconnect_2:VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, x_coordinate:reset_n, y_coordinate:reset_n]
	wire          rst_controller_reset_out_reset_req;                                   // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire          arm_a9_hps_h2f_reset_reset;                                           // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire          system_pll_reset_source_reset;                                        // System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> VGA_Subsystem:sys_reset_reset_n
	wire          rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                         //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                        //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                       //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                     //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),      //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),        //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),        //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),        //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),        //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),        //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),        //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),         //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),      //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),      //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),      //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),        //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),        //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),        //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),          //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),          //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),          //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),          //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),          //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),          //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),          //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),           //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),           //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),          //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),           //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),           //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),           //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),           //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),           //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),           //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),           //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),           //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),           //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),           //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),          //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),          //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),          //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),          //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),         //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),        //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),        //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),         //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),          //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),          //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),          //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),          //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),          //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),          //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),       //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),       //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),       //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),       //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),       //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),       //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),       //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),       //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID                 (arm_a9_hps_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR               (arm_a9_hps_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN                (arm_a9_hps_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE               (arm_a9_hps_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST              (arm_a9_hps_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK               (arm_a9_hps_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE              (arm_a9_hps_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT               (arm_a9_hps_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID              (arm_a9_hps_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY              (arm_a9_hps_h2f_axi_master_awready),    //                  .awready
		.h2f_WID                  (arm_a9_hps_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA                (arm_a9_hps_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB                (arm_a9_hps_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST                (arm_a9_hps_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID               (arm_a9_hps_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY               (arm_a9_hps_h2f_axi_master_wready),     //                  .wready
		.h2f_BID                  (arm_a9_hps_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP                (arm_a9_hps_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID               (arm_a9_hps_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY               (arm_a9_hps_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID                 (arm_a9_hps_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR               (arm_a9_hps_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN                (arm_a9_hps_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE               (arm_a9_hps_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST              (arm_a9_hps_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK               (arm_a9_hps_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE              (arm_a9_hps_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT               (arm_a9_hps_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID              (arm_a9_hps_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY              (arm_a9_hps_h2f_axi_master_arready),    //                  .arready
		.h2f_RID                  (arm_a9_hps_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA                (arm_a9_hps_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP                (arm_a9_hps_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST                (arm_a9_hps_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID               (arm_a9_hps_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY               (arm_a9_hps_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),               //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                     //                  .awaddr
		.f2h_AWLEN                (),                                     //                  .awlen
		.f2h_AWSIZE               (),                                     //                  .awsize
		.f2h_AWBURST              (),                                     //                  .awburst
		.f2h_AWLOCK               (),                                     //                  .awlock
		.f2h_AWCACHE              (),                                     //                  .awcache
		.f2h_AWPROT               (),                                     //                  .awprot
		.f2h_AWVALID              (),                                     //                  .awvalid
		.f2h_AWREADY              (),                                     //                  .awready
		.f2h_AWUSER               (),                                     //                  .awuser
		.f2h_WID                  (),                                     //                  .wid
		.f2h_WDATA                (),                                     //                  .wdata
		.f2h_WSTRB                (),                                     //                  .wstrb
		.f2h_WLAST                (),                                     //                  .wlast
		.f2h_WVALID               (),                                     //                  .wvalid
		.f2h_WREADY               (),                                     //                  .wready
		.f2h_BID                  (),                                     //                  .bid
		.f2h_BRESP                (),                                     //                  .bresp
		.f2h_BVALID               (),                                     //                  .bvalid
		.f2h_BREADY               (),                                     //                  .bready
		.f2h_ARID                 (),                                     //                  .arid
		.f2h_ARADDR               (),                                     //                  .araddr
		.f2h_ARLEN                (),                                     //                  .arlen
		.f2h_ARSIZE               (),                                     //                  .arsize
		.f2h_ARBURST              (),                                     //                  .arburst
		.f2h_ARLOCK               (),                                     //                  .arlock
		.f2h_ARCACHE              (),                                     //                  .arcache
		.f2h_ARPROT               (),                                     //                  .arprot
		.f2h_ARVALID              (),                                     //                  .arvalid
		.f2h_ARREADY              (),                                     //                  .arready
		.f2h_ARUSER               (),                                     //                  .aruser
		.f2h_RID                  (),                                     //                  .rid
		.f2h_RDATA                (),                                     //                  .rdata
		.f2h_RRESP                (),                                     //                  .rresp
		.f2h_RLAST                (),                                     //                  .rlast
		.f2h_RVALID               (),                                     //                  .rvalid
		.f2h_RREADY               (),                                     //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	Computer_System_AV_Config av_config (
		.clk         (system_pll_sys_clk_clk),                                         //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_1_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_1_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_1_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_1_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_1_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_1_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                  //                       .export
	);

	Computer_System_Onchip_SRAM onchip_sram (
		.address     (),                                            //     s1.address
		.clken       (),                                            //       .clken
		.chipselect  (),                                            //       .chipselect
		.write       (),                                            //       .write
		.readdata    (),                                            //       .readdata
		.writedata   (),                                            //       .writedata
		.address2    (mm_interconnect_0_onchip_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_sram_s2_writedata),  //       .writedata
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) pixel_dma_addr_translation (
		.clk                (system_pll_sys_clk_clk),                                         //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                 //  reset.reset
		.slave_address      (mm_interconnect_1_pixel_dma_addr_translation_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_1_pixel_dma_addr_translation_slave_read),        //       .read
		.slave_write        (mm_interconnect_1_pixel_dma_addr_translation_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_1_pixel_dma_addr_translation_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_1_pixel_dma_addr_translation_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest), //       .waitrequest
		.master_readdata    (pixel_dma_addr_translation_master_readdata),                     // master.readdata
		.master_waitrequest (pixel_dma_addr_translation_master_waitrequest),                  //       .waitrequest
		.master_address     (pixel_dma_addr_translation_master_address),                      //       .address
		.master_byteenable  (pixel_dma_addr_translation_master_byteenable),                   //       .byteenable
		.master_read        (pixel_dma_addr_translation_master_read),                         //       .read
		.master_write       (pixel_dma_addr_translation_master_write),                        //       .write
		.master_writedata   (pixel_dma_addr_translation_master_writedata)                     //       .writedata
	);

	Computer_System_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_VGA_Subsystem vga_subsystem (
		.char_buffer_control_slave_address    (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_chipselect (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect), //                          .chipselect
		.char_buffer_control_slave_read       (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_byteenable         (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),         //         char_buffer_slave.byteenable
		.char_buffer_slave_chipselect         (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_read               (mm_interconnect_0_vga_subsystem_char_buffer_slave_read),               //                          .read
		.char_buffer_slave_write              (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_writedata          (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_readdata           (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_waitrequest        (mm_interconnect_0_vga_subsystem_char_buffer_slave_waitrequest),        //                          .waitrequest
		.char_buffer_slave_address            (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),            //                          .address
		.pixel_dma_control_slave_address      (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_readdata),     //                          .readdata
		.pixel_dma_master_readdatavalid       (vga_subsystem_pixel_dma_master_readdatavalid),                         //          pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest         (vga_subsystem_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_address             (vga_subsystem_pixel_dma_master_address),                               //                          .address
		.pixel_dma_master_lock                (vga_subsystem_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vga_subsystem_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vga_subsystem_pixel_dma_master_readdata),                              //                          .readdata
		.sys_clk_clk                          (system_pll_sys_clk_clk),                                               //                   sys_clk.clk
		.sys_reset_reset_n                    (~rst_controller_001_reset_out_reset),                                  //                 sys_reset.reset_n
		.vga_CLK                              (vga_CLK),                                                              //                       vga.CLK
		.vga_HS                               (vga_HS),                                                               //                          .HS
		.vga_VS                               (vga_VS),                                                               //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                            //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                             //                          .SYNC
		.vga_R                                (vga_R),                                                                //                          .R
		.vga_G                                (vga_G),                                                                //                          .G
		.vga_B                                (vga_B),                                                                //                          .B
		.vga_pll_ref_clk_clk                  (vga_pll_ref_clk_clk),                                                  //           vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset              (vga_pll_ref_reset_reset)                                               //         vga_pll_ref_reset.reset
	);

	Computer_System_x_coordinate x_coordinate (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_x_coordinate_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_x_coordinate_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_x_coordinate_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_x_coordinate_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_x_coordinate_s1_readdata),   //                    .readdata
		.out_port   (x_coordinate_external_connection_export)       // external_connection.export
	);

	Computer_System_x_coordinate y_coordinate (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_y_coordinate_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_y_coordinate_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_y_coordinate_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_y_coordinate_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_y_coordinate_s1_readdata),   //                    .readdata
		.out_port   (y_coordinate_external_connection_export)       // external_connection.export
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),                                //                                       ARM_A9_HPS_h2f_axi_master.awid
		.ARM_A9_HPS_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),                              //                                                                .awaddr
		.ARM_A9_HPS_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),                               //                                                                .awlen
		.ARM_A9_HPS_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),                              //                                                                .awsize
		.ARM_A9_HPS_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),                             //                                                                .awburst
		.ARM_A9_HPS_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),                              //                                                                .awlock
		.ARM_A9_HPS_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),                             //                                                                .awcache
		.ARM_A9_HPS_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),                              //                                                                .awprot
		.ARM_A9_HPS_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),                             //                                                                .awvalid
		.ARM_A9_HPS_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),                             //                                                                .awready
		.ARM_A9_HPS_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),                                 //                                                                .wid
		.ARM_A9_HPS_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),                               //                                                                .wdata
		.ARM_A9_HPS_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),                               //                                                                .wstrb
		.ARM_A9_HPS_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),                               //                                                                .wlast
		.ARM_A9_HPS_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),                              //                                                                .wvalid
		.ARM_A9_HPS_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),                              //                                                                .wready
		.ARM_A9_HPS_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),                                 //                                                                .bid
		.ARM_A9_HPS_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),                               //                                                                .bresp
		.ARM_A9_HPS_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),                              //                                                                .bvalid
		.ARM_A9_HPS_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),                              //                                                                .bready
		.ARM_A9_HPS_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),                                //                                                                .arid
		.ARM_A9_HPS_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),                              //                                                                .araddr
		.ARM_A9_HPS_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),                               //                                                                .arlen
		.ARM_A9_HPS_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),                              //                                                                .arsize
		.ARM_A9_HPS_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),                             //                                                                .arburst
		.ARM_A9_HPS_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),                              //                                                                .arlock
		.ARM_A9_HPS_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),                             //                                                                .arcache
		.ARM_A9_HPS_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),                              //                                                                .arprot
		.ARM_A9_HPS_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),                             //                                                                .arvalid
		.ARM_A9_HPS_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),                             //                                                                .arready
		.ARM_A9_HPS_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),                                 //                                                                .rid
		.ARM_A9_HPS_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),                               //                                                                .rdata
		.ARM_A9_HPS_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),                               //                                                                .rresp
		.ARM_A9_HPS_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),                               //                                                                .rlast
		.ARM_A9_HPS_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),                              //                                                                .rvalid
		.ARM_A9_HPS_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),                              //                                                                .rready
		.System_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                                        //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                            // ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.SDRAM_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                                //                               SDRAM_reset_reset_bridge_in_reset.reset
		.VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                                //                   VGA_Subsystem_sys_reset_reset_bridge_in_reset.reset
		.VGA_Subsystem_pixel_dma_master_address                                (vga_subsystem_pixel_dma_master_address),                        //                                  VGA_Subsystem_pixel_dma_master.address
		.VGA_Subsystem_pixel_dma_master_waitrequest                            (vga_subsystem_pixel_dma_master_waitrequest),                    //                                                                .waitrequest
		.VGA_Subsystem_pixel_dma_master_read                                   (vga_subsystem_pixel_dma_master_read),                           //                                                                .read
		.VGA_Subsystem_pixel_dma_master_readdata                               (vga_subsystem_pixel_dma_master_readdata),                       //                                                                .readdata
		.VGA_Subsystem_pixel_dma_master_readdatavalid                          (vga_subsystem_pixel_dma_master_readdatavalid),                  //                                                                .readdatavalid
		.VGA_Subsystem_pixel_dma_master_lock                                   (vga_subsystem_pixel_dma_master_lock),                           //                                                                .lock
		.Onchip_SRAM_s2_address                                                (mm_interconnect_0_onchip_sram_s2_address),                      //                                                  Onchip_SRAM_s2.address
		.Onchip_SRAM_s2_write                                                  (mm_interconnect_0_onchip_sram_s2_write),                        //                                                                .write
		.Onchip_SRAM_s2_readdata                                               (mm_interconnect_0_onchip_sram_s2_readdata),                     //                                                                .readdata
		.Onchip_SRAM_s2_writedata                                              (mm_interconnect_0_onchip_sram_s2_writedata),                    //                                                                .writedata
		.Onchip_SRAM_s2_chipselect                                             (mm_interconnect_0_onchip_sram_s2_chipselect),                   //                                                                .chipselect
		.Onchip_SRAM_s2_clken                                                  (mm_interconnect_0_onchip_sram_s2_clken),                        //                                                                .clken
		.SDRAM_s1_address                                                      (mm_interconnect_0_sdram_s1_address),                            //                                                        SDRAM_s1.address
		.SDRAM_s1_write                                                        (mm_interconnect_0_sdram_s1_write),                              //                                                                .write
		.SDRAM_s1_read                                                         (mm_interconnect_0_sdram_s1_read),                               //                                                                .read
		.SDRAM_s1_readdata                                                     (mm_interconnect_0_sdram_s1_readdata),                           //                                                                .readdata
		.SDRAM_s1_writedata                                                    (mm_interconnect_0_sdram_s1_writedata),                          //                                                                .writedata
		.SDRAM_s1_byteenable                                                   (mm_interconnect_0_sdram_s1_byteenable),                         //                                                                .byteenable
		.SDRAM_s1_readdatavalid                                                (mm_interconnect_0_sdram_s1_readdatavalid),                      //                                                                .readdatavalid
		.SDRAM_s1_waitrequest                                                  (mm_interconnect_0_sdram_s1_waitrequest),                        //                                                                .waitrequest
		.SDRAM_s1_chipselect                                                   (mm_interconnect_0_sdram_s1_chipselect),                         //                                                                .chipselect
		.VGA_Subsystem_char_buffer_slave_address                               (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),     //                                 VGA_Subsystem_char_buffer_slave.address
		.VGA_Subsystem_char_buffer_slave_write                                 (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),       //                                                                .write
		.VGA_Subsystem_char_buffer_slave_read                                  (mm_interconnect_0_vga_subsystem_char_buffer_slave_read),        //                                                                .read
		.VGA_Subsystem_char_buffer_slave_readdata                              (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),    //                                                                .readdata
		.VGA_Subsystem_char_buffer_slave_writedata                             (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),   //                                                                .writedata
		.VGA_Subsystem_char_buffer_slave_byteenable                            (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),  //                                                                .byteenable
		.VGA_Subsystem_char_buffer_slave_waitrequest                           (mm_interconnect_0_vga_subsystem_char_buffer_slave_waitrequest), //                                                                .waitrequest
		.VGA_Subsystem_char_buffer_slave_chipselect                            (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect)   //                                                                .chipselect
	);

	Computer_System_mm_interconnect_1 mm_interconnect_1 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                                    //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                                  //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                                   //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                                  //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                                 //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                                  //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                                 //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                                  //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                                 //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                                 //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                                     //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                                   //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                                   //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                                   //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                                  //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                                  //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                                     //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                                   //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                                  //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                                  //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                                    //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                                  //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                                   //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                                  //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                                 //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                                  //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                                 //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                                  //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                                 //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                                 //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                                     //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                                   //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                                   //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                                   //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                                  //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                                  //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                               //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                   // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.AV_Config_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                       //                              AV_Config_reset_reset_bridge_in_reset.reset
		.VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                                       //                      VGA_Subsystem_sys_reset_reset_bridge_in_reset.reset
		.AV_Config_avalon_av_config_slave_address                                 (mm_interconnect_1_av_config_avalon_av_config_slave_address),           //                                   AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                                   (mm_interconnect_1_av_config_avalon_av_config_slave_write),             //                                                                   .write
		.AV_Config_avalon_av_config_slave_read                                    (mm_interconnect_1_av_config_avalon_av_config_slave_read),              //                                                                   .read
		.AV_Config_avalon_av_config_slave_readdata                                (mm_interconnect_1_av_config_avalon_av_config_slave_readdata),          //                                                                   .readdata
		.AV_Config_avalon_av_config_slave_writedata                               (mm_interconnect_1_av_config_avalon_av_config_slave_writedata),         //                                                                   .writedata
		.AV_Config_avalon_av_config_slave_byteenable                              (mm_interconnect_1_av_config_avalon_av_config_slave_byteenable),        //                                                                   .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest                             (mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest),       //                                                                   .waitrequest
		.Pixel_DMA_Addr_Translation_slave_address                                 (mm_interconnect_1_pixel_dma_addr_translation_slave_address),           //                                   Pixel_DMA_Addr_Translation_slave.address
		.Pixel_DMA_Addr_Translation_slave_write                                   (mm_interconnect_1_pixel_dma_addr_translation_slave_write),             //                                                                   .write
		.Pixel_DMA_Addr_Translation_slave_read                                    (mm_interconnect_1_pixel_dma_addr_translation_slave_read),              //                                                                   .read
		.Pixel_DMA_Addr_Translation_slave_readdata                                (mm_interconnect_1_pixel_dma_addr_translation_slave_readdata),          //                                                                   .readdata
		.Pixel_DMA_Addr_Translation_slave_writedata                               (mm_interconnect_1_pixel_dma_addr_translation_slave_writedata),         //                                                                   .writedata
		.Pixel_DMA_Addr_Translation_slave_byteenable                              (mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable),        //                                                                   .byteenable
		.Pixel_DMA_Addr_Translation_slave_waitrequest                             (mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest),       //                                                                   .waitrequest
		.VGA_Subsystem_char_buffer_control_slave_address                          (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address),    //                            VGA_Subsystem_char_buffer_control_slave.address
		.VGA_Subsystem_char_buffer_control_slave_write                            (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write),      //                                                                   .write
		.VGA_Subsystem_char_buffer_control_slave_read                             (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read),       //                                                                   .read
		.VGA_Subsystem_char_buffer_control_slave_readdata                         (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata),   //                                                                   .readdata
		.VGA_Subsystem_char_buffer_control_slave_writedata                        (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata),  //                                                                   .writedata
		.VGA_Subsystem_char_buffer_control_slave_byteenable                       (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable), //                                                                   .byteenable
		.VGA_Subsystem_char_buffer_control_slave_chipselect                       (mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect), //                                                                   .chipselect
		.x_coordinate_s1_address                                                  (mm_interconnect_1_x_coordinate_s1_address),                            //                                                    x_coordinate_s1.address
		.x_coordinate_s1_write                                                    (mm_interconnect_1_x_coordinate_s1_write),                              //                                                                   .write
		.x_coordinate_s1_readdata                                                 (mm_interconnect_1_x_coordinate_s1_readdata),                           //                                                                   .readdata
		.x_coordinate_s1_writedata                                                (mm_interconnect_1_x_coordinate_s1_writedata),                          //                                                                   .writedata
		.x_coordinate_s1_chipselect                                               (mm_interconnect_1_x_coordinate_s1_chipselect),                         //                                                                   .chipselect
		.y_coordinate_s1_address                                                  (mm_interconnect_1_y_coordinate_s1_address),                            //                                                    y_coordinate_s1.address
		.y_coordinate_s1_write                                                    (mm_interconnect_1_y_coordinate_s1_write),                              //                                                                   .write
		.y_coordinate_s1_readdata                                                 (mm_interconnect_1_y_coordinate_s1_readdata),                           //                                                                   .readdata
		.y_coordinate_s1_writedata                                                (mm_interconnect_1_y_coordinate_s1_writedata),                          //                                                                   .writedata
		.y_coordinate_s1_chipselect                                               (mm_interconnect_1_y_coordinate_s1_chipselect)                          //                                                                   .chipselect
	);

	Computer_System_mm_interconnect_2 mm_interconnect_2 (
		.System_PLL_sys_clk_clk                                       (system_pll_sys_clk_clk),                                             //                                     System_PLL_sys_clk.clk
		.Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset.reset
		.VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                     //          VGA_Subsystem_sys_reset_reset_bridge_in_reset.reset
		.Pixel_DMA_Addr_Translation_master_address                    (pixel_dma_addr_translation_master_address),                          //                      Pixel_DMA_Addr_Translation_master.address
		.Pixel_DMA_Addr_Translation_master_waitrequest                (pixel_dma_addr_translation_master_waitrequest),                      //                                                       .waitrequest
		.Pixel_DMA_Addr_Translation_master_byteenable                 (pixel_dma_addr_translation_master_byteenable),                       //                                                       .byteenable
		.Pixel_DMA_Addr_Translation_master_read                       (pixel_dma_addr_translation_master_read),                             //                                                       .read
		.Pixel_DMA_Addr_Translation_master_readdata                   (pixel_dma_addr_translation_master_readdata),                         //                                                       .readdata
		.Pixel_DMA_Addr_Translation_master_write                      (pixel_dma_addr_translation_master_write),                            //                                                       .write
		.Pixel_DMA_Addr_Translation_master_writedata                  (pixel_dma_addr_translation_master_writedata),                        //                                                       .writedata
		.VGA_Subsystem_pixel_dma_control_slave_address                (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_address),    //                  VGA_Subsystem_pixel_dma_control_slave.address
		.VGA_Subsystem_pixel_dma_control_slave_write                  (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_write),      //                                                       .write
		.VGA_Subsystem_pixel_dma_control_slave_read                   (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_read),       //                                                       .read
		.VGA_Subsystem_pixel_dma_control_slave_readdata               (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_readdata),   //                                                       .readdata
		.VGA_Subsystem_pixel_dma_control_slave_writedata              (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_writedata),  //                                                       .writedata
		.VGA_Subsystem_pixel_dma_control_slave_byteenable             (mm_interconnect_2_vga_subsystem_pixel_dma_control_slave_byteenable)  //                                                       .byteenable
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
